SIGNAL tx_buffer      : tx_array :=
(

	"010000000000001000100011010001000000000000000111",
	"010000000000001000100011100001000000000000000000",
	"010000000000001000100011010001000100000000000111",
	"010000000000001000100011100001000000000000010000",
	"010000000000010000100011010001000000000000000111",
	"010000000000010000100011100001000000000000000000",
	"010000000000010000100011010001000100000000000111",
	"010000000000010000100011100001000000000000010000",
	"010000000000011000100011010001000000000000000111",
	"010000000000011000100011100001000000000000000000",
	"010000000000011000100011010001000100000000000111",
	"010000000000011000100011100001000000000000010000",
	"010000000000100000100011010001000000000000000111",
	"010000000000100000100011100001000000000000000000",
	"010000000000100000100011010001000100000000000111",
	"010000000000100000100011100001000000000000010000",
	"010000000000101000100011010001000000000000000111",
	"010000000000101000100011100001000000000000000000",
	"010000000000101000100011010001000100000000000111",
	"010000000000101000100011100001000000000000010000",
	"010000000000001000100011010001000000000000000111",
	"010000000000001000100011100001000000000000111100",
	"010000000000001000100011010001000100000000000111",
	"010000000000001000100011100001000000000000000000",
	"010000000000010000100011010001000000000000000111",
	"010000000000010000100011100001000000000000111100",
	"010000000000010000100011010001000100000000000111",
	"010000000000010000100011100001000000000000000000",
	"010000000000011000100011010001000000000000000111",
	"010000000000011000100011100001000000000000111100",
	"010000000000011000100011010001000100000000000111",
	"010000000000011000100011100001000000000000000000",
	"010000000000100000100011010001000000000000000111",
	"010000000000100000100011100001000000000000111100",
	"010000000000100000100011010001000100000000000111",
	"010000000000100000100011100001000000000000000000",
	"010000000000101000100011010001000000000000000111",
	"010000000000101000100011100001000000000000111100",
	"010000000000101000100011010001000100000000000111",
	"010000000000101000100011100001000000000000000000",

);